`timescale 1 ps / 1 ps

module design_1_wrapper
   (clk_0);
  input clk_0;

  wire clk_0;

  design_1 design_1_i
       (.clk_0(clk_0));
endmodule
